library ieee;
use ieee.std_logic_1164.all; 
use work.all;

entity multimedia_alu_tb is
end entity;

architecture testbench of multimedia_alu_tb is 

signal rs1, rs2, rs3, rd: std_logic_vector(127 downto 0);
signal rd_add, rd_addr : std_logic_vector(4 downto 0);
signal opcode: std_logic_vector(7 downto 0);
signal instr: std_logic_vector(1 downto 0);	 
signal load_index : std_logic_vector (2 downto 0);	
signal imm : std_logic_vector (15 downto 0);

component multimedia_alu
    port (										 
        rs1 : in std_logic_vector (127 downto 0);
		rs2 : in std_logic_vector (127 downto 0);
		rs3 : in std_logic_vector (127 downto 0); 
		opcode : in std_logic_vector (7 downto 0); 
		load_index : in std_logic_vector (2 downto 0);
		imm : in std_logic_vector (15 downto 0);
		instr : in std_logic_vector (1 downto 0);	 
		rd : out std_logic_vector (127 downto 0)
    );
end component;

begin
    uut: entity multimedia_alu
        port map (
            rs1 => rs1,
            rs2 => rs2,
            rs3 => rs3,	 	   
            opcode => opcode,
			load_index => load_index,
			imm => imm,
            instr => instr,
            rd => rd
        );

    stimulus: process
    begin	 
		
		wait for 10ns;
		
		rs1 <= x"00000000000000000000000000000032";
        rs2 <= x"00000000FFFF00000000000000000003";
        rs3 <= x"00000000FFFF00000000000000000064";	
		instr <= "10";
		opcode <= "-----000";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----001";
        wait for 20 ns;
		report "rd = " & to_string(rd);	   
		
		
		
		wait for 10ns;	 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----010";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----011";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----100";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "00000000000000000000000000000000" & "00000000000000000000000000001010" & "00000000000000000000000000000000" & "00000000000000000000000000101000";
        rs2 <= "00000000000000000000000000000000" & "00000000000000000000000000000001" & "00000000000000000000000000000000" & "00000000000000000000000000000100";
        rs3 <= "00000000000000000000000000000000" & "00000000000000000000000000000101" & "00000000000000000000000000000000" & "00000000000000000000000000000101";	
		instr <= "10";
		opcode <= "-----110";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----111";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----000";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----001";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----010";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----011";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----100";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "10";
		opcode <= "-----110";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0001";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "00000000000000000000000000000000" & "00000000000000000000000000000001" & "00000000000000000000000000000000" & "00000000000000000000000000000100";
        rs2 <= "00000000000000000000000000000000" & "00000000000000000000000000000101" & "00000000000000000000000000000000" & "00000000000000000000000000000101";	
		instr <= "11";
		opcode <= "----0010";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0011";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0100";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0110";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----0111";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "---01000";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	   
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1001";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "10000000000000000000000000000000000000001000000000000000000000000000000000000000000000011000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1010";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "10000000000000000000000000000000000000001000000000000000000000000000000000000000000000011000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000010000000000000000000000000000000000000000000011000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1011";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1100";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;	
		
		rs1 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1110";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		rs1 <= "00001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
        rs2 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100";
        rs3 <= "10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";	
		instr <= "11";
		opcode <= "----1111";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		
		rs1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        instr <= "0-";
		load_index <= "000";   
		imm <= "0001101110110101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns; 
		
		rs1 <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101110110101";
        instr <= "0-";
		load_index <= "111";   
		imm <= "0001101110110101";
        wait for 20 ns;
		report "rd = " & to_string(rd);	  
		
		wait for 10ns;
		
		
		wait;
		
		wait;
		
	end process;
end testbench;
